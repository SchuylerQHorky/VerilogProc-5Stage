/**********************************************************8
Instruction Fetch, takes in the next instruction ,determines 
which kind of instruction it is and then breaks it apart into
its constituent pieces to pass to the rest of the processor


************************************************************/

module inst_fetch (instructions, br_taken, zero, overflow, negative, condAddr) begin




end module